// module ysyx_23060061_UART (
// 	input clk,
// 	input rst, // low activate
//
// 	input [31:0] araddr,
// 	input arvalid,
// 	output reg arready,
//
// 	output reg [31:0] rdata,
// 	output reg [1:0] rresp,
// 	output reg rvalid,
// 	input rready,
//
// 	input [31:0] awaddr,
// 	input awvalid,
// 	output reg awready,
//
// 	input [31:0] wdata,
// 	input [3:0] wstrb,
// 	input wvalid,
// 	output reg wready,
//
// 	output reg [1:0] bresp,
// 	output reg bvalid,
// 	input bready
// );
// 	// FSM
// 	reg [2:0] state;
// 	localparam   = ;	
// endmodule