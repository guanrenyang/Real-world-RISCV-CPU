// module ysyx