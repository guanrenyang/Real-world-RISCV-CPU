// module ysyx_23060061_WB(
// 	input clk,
// 	input rst,
//
// 	input [31:0] memDataR,
// 	input [31:0] aluOut,
// 	input [31:0] snpc,
// 	input [31:0] dnpc,
// 	input [31:0] csrReadData;
//
// );
// endmodule