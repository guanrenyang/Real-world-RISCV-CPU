module ysyx_23060061_Decoder (
  input [6:0] opcode,
  input [2:0] funct3
);
  

endmodule
