module ysyx_23060061_BranchComp(
	input [31:0] rdata1,
	input [31:0] rdata2,
	input BrUn, // branch unsigned
	output BrEq,
	output BrLt
);

endmodule